*** inverter ***
.subckt inv Vin Vout VDD GND
MnMos Vout Vin GND GND n_18 W=0.5u L=0.18u
MpMos Vout Vin VDD VDD p_18 W=1u L=0.18u
.ends

*** nand ***
.subckt nand A B out_2 VDD GND
MnMos1 out_2 A net1 GND n_18 W=0.5u L=0.18u
MnMos2 net1 B GND GND n_18 W=0.5u L=0.18u
MpMos1 out_2 A VDD VDD p_18 W=1u L=0.18u
MpMos2 out_2 B VDD VDD p_18 W=1u L=0.18u
.ends

*** nor ***
.subckt nor C D out_3 VDD GND
MnMos1 out_3 C GND GND n_18 W=0.5u L=0.18u
MnMos2 out_3 D GND GND n_18 W=0.5u L=0.18u
MpMos1 net1 C VDD VDD p_18 W=1u L=0.18u
MpMos2 out_3 D net1 VDD p_18 W=1u L=0.18u
.ends
