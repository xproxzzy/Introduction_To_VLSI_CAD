.INC 'fulladder.spi'
*** RCA ***
.subckt RCA A0 B0 C0 A1 B1 A2 B2 A3 B3 C4 S0 S1 S2 S3 VDD GND
Xfulladder0 A0 B0 C0 S0 C1 VDD GND fulladder
Xfulladder1 A1 B1 C1 S1 C2 VDD GND fulladder
Xfulladder2 A2 B2 C2 S2 C3 VDD GND fulladder
Xfulladder3 A3 B3 C3 S3 C4 VDD GND fulladder
.ends
