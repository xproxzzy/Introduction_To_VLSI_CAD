*** halfadder ***
.subckt halfadder X Y S C VDD GND
MnMos5 neg_X X GND GND n_18 W=0.5u L=0.18u
MpMos5 neg_X X VDD VDD p_18 W=1u L=0.18u
MnMos6 neg_Y Y GND GND n_18 W=0.5u L=0.18u
MpMos6 neg_Y Y VDD VDD p_18 W=1u L=0.18u
MpMos1 net1 neg_X VDD VDD p_18 W=1u L=0.18u
MpMos2 S Y net1 VDD p_18 W=1u L=0.18u
MpMos3 net2 X VDD VDD p_18 W=1u L=0.18u
MpMos4 S neg_Y net2 VDD p_18 W=1u L=0.18u
MnMos1 S neg_Y net3 GND n_18 W=0.5u L=0.18u
MnMos2 net3 Y GND GND n_18 W=0.5u L=0.18u
MnMos3 S X net3 GND n_18 W=0.5u L=0.18u
MnMos4 net3 neg_X GND GND n_18 W=0.5u L=0.18u
MnMos7 net5 X net4 GND n_18 W=0.5u L=0.18u
MnMos8 net4 Y GND GND n_18 W=0.5u L=0.18u
MpMos7 net5 X VDD VDD p_18 W=1u L=0.18u
MpMos8 net5 Y VDD VDD p_18 W=1u L=0.18u
MnMos9 C net5 GND GND n_18 W=0.5u L=0.18u
MpMos9 C net5 VDD VDD p_18 W=1u L=0.18u
.ends
